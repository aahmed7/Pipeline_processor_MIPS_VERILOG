module ALUsub(func,ALUOp,ALUCtrl);
	input [5:0]func;
	input [1:0]ALUOp;
	output [3:0]ALUCtrl